LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY dec4to16 IS
	PORT (w  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0) ;
			En : IN  STD_LOGIC ;
			Y:  OUT STD_LOGIC_VECTOR(15 downto 0))  ;
		
END ENTITY ;

ARCHITECTURE Behavior OF dec4to16 IS
	SIGNAL Enw : STD_LOGIC_VECTOR(4 DOWNTO 0) ;
BEGIN
	Enw <= En & w ;
	WITH Enw SELECT
	Y <=    "1000000000000000" WHEN "10000", -- 0
           "0100000000000000" WHEN "10001", -- 1
           "0010000000000000" WHEN "10010", -- 2
           "0001000000000000" WHEN "10011", -- 3
           "0000100000000000" WHEN "10100", -- 4
           "0000010000000000" WHEN "10101", -- 5
           "0000001000000000" WHEN "10110", -- 6
			  "0000000100000000" WHEN "10111", -- 7
           "0000000010000000" WHEN "11000", -- 8
           "0000000001000000" WHEN "11001", -- 9
           "0000000000100000" WHEN "11010", -- 10
           "0000000000010000" WHEN "11011", -- 11
           "0000000000001000" WHEN "11100", -- 12
           "0000000000000100" WHEN "11101", -- 13
           "0000000000000010" WHEN "11110", -- 14
           "0000000000000001" WHEN "11111", -- 15
           "0000000000000000" WHEN OTHERS;  -- Dont care
		
END Behavior ;