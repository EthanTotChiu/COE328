library verilog;
use verilog.vl_types.all;
entity Lab6_problem3_vlg_vec_tst is
end Lab6_problem3_vlg_vec_tst;
